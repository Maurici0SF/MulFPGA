library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use ieee.std_logic_unsigned.all;
entity W is
	port (Spike,CLK: 	in STD_LOGIC;
			Num:		out STD_LOGIC_VECTOR(3 downto 0));
end W;

architecture behav of W is
	
begin
	
end behav;